library IEEE;
use IEEE.std_logic_1164.all;

entity Decoder6t64 is
    port(input : in std_logic_vector(5 downto 0);
        output : out std_logic_vector(63 downto 0));
end Decoder6t64;

architecture dataflow of Decoder6t64 is
begin
    with input select output <= 
        x"0000000000000001" when "000000",
        x"0000000000000002" when "000001",
        x"0000000000000004" when "000010",
        x"0000000000000008" when "000011",
        x"0000000000000010" when "000100",
        x"0000000000000020" when "000101",
        x"0000000000000040" when "000110",
        x"0000000000000080" when "000111",
        x"0000000000000100" when "001000",
        x"0000000000000200" when "001001",
        x"0000000000000400" when "001010",
        x"0000000000000800" when "001011",
        x"0000000000001000" when "001100",
        x"0000000000002000" when "001101",
        x"0000000000004000" when "001110",
        x"0000000000008000" when "001111",
        x"0000000000010000" when "010000",
        x"0000000000020000" when "010001",
        x"0000000000040000" when "010010",
        x"0000000000080000" when "010011",
        x"0000000000100000" when "010100",
        x"0000000000200000" when "010101",
        x"0000000000400000" when "010110",
        x"0000000000800000" when "010111",
        x"0000000001000000" when "011000",
        x"0000000002000000" when "011001",
        x"0000000004000000" when "011010",
        x"0000000008000000" when "011011",
        x"0000000010000000" when "011100",
        x"0000000020000000" when "011101",
        x"0000000040000000" when "011110",
        x"0000000080000000" when "011111",
        x"0000000100000000" when "100000",
        x"0000000200000000" when "100001",
        x"0000000400000000" when "100010",
        x"0000000800000000" when "100011",
        x"0000001000000000" when "100100",
        x"0000002000000000" when "100101",
        x"0000004000000000" when "100110",
        x"0000008000000000" when "100111",
        x"0000010000000000" when "101000",
        x"0000020000000000" when "101001",
        x"0000040000000000" when "101010",
        x"0000080000000000" when "101011",
        x"0000100000000000" when "101100",
        x"0000200000000000" when "101101",
        x"0000400000000000" when "101110",
        x"0000800000000000" when "101111",
        x"0001000000000000" when "110000",
        x"0002000000000000" when "110001",
        x"0004000000000000" when "110010",
        x"0008000000000000" when "110011",
        x"0010000000000000" when "110100",
        x"0020000000000000" when "110101",
        x"0040000000000000" when "110110",
        x"0080000000000000" when "110111",
        x"0100000000000000" when "111000",
        x"0200000000000000" when "111001",
        x"0400000000000000" when "111010",
        x"0800000000000000" when "111011",
        x"1000000000000000" when "111100",
        x"2000000000000000" when "111101",
        x"4000000000000000" when "111110",
        x"8000000000000000" when "111111",
        x"0000000000000000" when others;
end dataflow;